module gt10(
	input [3:0]a,
	output b
);
assign b = a > 10 ? 1 : 0;
endmodule
