module reg_fl_tb;
reg clk, rst_b,[7:0]wr_data; reg [1:0]wr_addr; reg wr_l,[1:0]rd_addr; reg rd_l;
wire [7:0]rd_data;
