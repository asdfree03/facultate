module comparator(
	input [1:0]x, 
	input [1:0]y,
	output eq,le,gt
);
	assign eq = ((~x[1]) && (~x[0]) && (~y[1]) && (~y[0])) || ((~x[1]) && x[0] && (~y[1]) && y[0]) || (x[1] && x[0] && y[1] && y[0]) || (x[1] && (~x[0]) && y[1] && (~y[0]));
	assign le = ((~x[1]) && (~x[0]) && y[0]) || ((~x[0]) && y[1] && y[0]) || ((~x[1]) && y[1]);
	assign gt = (x[0] && (~y[1]) && (~y[0])) || (x[1] && x[0] && (~y[0])) || (x[1] && (~y[1]));
endmodule
